module example(
);
endmodule
